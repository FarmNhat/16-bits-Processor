module int_float(
);

endmodule